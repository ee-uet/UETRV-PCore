// Copyright 2023 University of Engineering and Technology Lahore.
// Licensed under the Apache License, Version 2.0, see LICENSE file for details.
// SPDX-License-Identifier: Apache-2.0
//
// Description:  A top level module for the 16 bit compressed instruction support.
//
// Author: Ateeb Tahir, DDRC, UET Lahore
// Date: 21.7.2023


